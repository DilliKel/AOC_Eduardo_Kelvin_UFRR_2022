-----------------------------------------------------------
-- COMPONENTE: BANCO DE REGISTRADORES
-- DESCRIÇÃO: 
--     ARMAZENA REGISTRADORES, PERMITINDO QUE NELES SEJAM
--     ESCRITOS E LIDOS DADOS
-----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BANCO_REGISTRADORES IS
    PORT(
        CLOCK,REG_WRITE     : IN STD_LOGIC;
        REG1_IN,REG2_IN     : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
        WRITE_DATA          : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        REG1_OUT,REG2_OUT  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END BANCO_REGISTRADORES;

ARCHITECTURE BEHAVIOR OF BANCO_REGISTRADORES IS
TYPE BANCO_DE_REGISTRADORES IS ARRAY(0 TO 3) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL MEM_BANCO_REG : BANCO_DE_REGISTRADORES;
BEGIN
    PROCESS(CLOCK,REG1_IN,REG2_IN,MEM_BANCO_REG)
    BEGIN
        IF RISING_EDGE(CLOCK) THEN
            IF (REG_WRITE = '1') THEN
                MEM_BANCO_REG(TO_INTEGER(UNSIGNED(REG1_IN))) <= WRITE_DATA;
            END IF;
        END IF;
        REG1_OUT <= MEM_BANCO_REG(TO_INTEGER(UNSIGNED(REG1_IN)));
        REG2_OUT <= MEM_BANCO_REG(TO_INTEGER(UNSIGNED(REG2_IN)));
    END PROCESS;
END;